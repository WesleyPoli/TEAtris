module teatris_memoria_mapas_dificil (
    input clock,                // Clock do sistema
    input [3:0] endereco,       // Endereço de memória (0-15)
    output reg [63:0] padrao     // Padrão de mapa para exibição
);

    // Memória ROM de padrões para mapas
    always @(posedge clock) begin
        case (endereco)
            
            4'd0: padrao <= {8'b000000_01,//8'b11_00_00_11,
                             8'b000000_11,//8'b11_01_01_11,
                             8'b001000_00,//8'b11_11_11_11,
                             8'b000100_00,//8'b11_00_00_11,
                             8'b110000_00,//8'b11_11_11_11,
                             8'b110000_00,//8'b11_00_00_11,
                             8'b000010_00,//8'b11_10_11_11,
                             8'b000011_00};//8'b11_00_00_11 //1

            4'd1: padrao <= {8'b00000010,
                             8'b00000010,
                             8'b00100000,
                             8'b01000000,
                             8'b00000010,
                             8'b00000110,
                             8'b0_11_00000,
                             8'b0_11_00000}; //4
            
            4'd2: padrao <= {8'b00000000,
                             8'b01100000,
                             8'b00001000,
                             8'b00001000,
                             8'b01100000,
                             8'b01000000,
                             8'b00000011,
                             8'b00000011}; //2 
                             
            4'd3: padrao <= {8'b00000001,
                             8'b00000010,
                             8'b00110000,
                             8'b00010000,
                             8'b00000000,
                             8'b00011000,
                             8'b10000000,
                             8'b11000000}; //3
                        
            4'd4: padrao <= {8'b01000000,
                             8'b11000000,
                             8'b00010000,
                             8'b00011000,
                             8'b01000000,
                             8'b00100000,
                             8'b00000010,
                             8'b00000010}; //2 

            4'd5: padrao <= {8'b00000011,
                             8'b00000001,
                             8'b00110000,
                             8'b00000000,
                             8'b00000011,
                             8'b00000011,
                             8'b00011000,
                             8'b00010000}; //4 
            
            4'd6: padrao <= {8'b00010000,
                             8'b00011000,
                             8'b01000000,
                             8'b00100000,
                             8'b00001000,
                             8'b00010000,
                             8'b00000110,
                             8'b00000010}; //3 
                             
            4'd7: padrao <= {8'b000_10_000,
                             8'b000_01_000,
                             8'b00100000,
                             8'b01100000,
                             8'b00001000,
                             8'b00001000,
                             8'b01100000,
                             8'b00100000}; //1 
                        
            4'd8: padrao <= {8'b00100000,
                             8'b01000000,
                             8'b00001100,
                             8'b00001000,
                             8'b01100000,
                             8'b00000000,
                             8'b00001000,
                             8'b00011000}; //4 

            4'd9: padrao <= {8'b00000001,
                             8'b00000011,
                             8'b10000000, 
                             8'b01000000, 
                             8'b00011000,
                             8'b00010000,
                             8'b00001000,
                             8'b00001100}; //3
            
            4'd10: padrao <= {8'b00001000,
                              8'b00010000,
                              8'b01000000,
                              8'b00100000,
                              8'b00000110,
                              8'b00000110,
                              8'b00110000,
                              8'b00100000}; //1 
                             
            4'd11: padrao <= {8'b00000001,
                              8'b00000011,
                              8'b00011000,
                              8'b00001000,
                              8'b11000000,
                              8'b11000000,
                              8'b00001000,
                              8'b00001100}; //2 
            4'd12: padrao <= {8'b00000001,
                              8'b00000011,
                              8'b10000000,
                              8'b01000000,
                              8'b00001100,
                              8'b00000000,
                              8'b01000000,
                              8'b01100000}; //3

            4'd13: padrao <= {8'b00011000,
                              8'b00011000,
                              8'b01000000,
                              8'b00100000,
                              8'b00000010,
                              8'b00000110,
                              8'b00100000,
                              8'b00110000}; //1 
            
            4'd14: padrao <= {8'b00000011,
                              8'b00000001,
                              8'b00010000,
                              8'b00010000,
                              8'b01000000,
                              8'b10000000,
                              8'b00001100,
                              8'b00001100}; //2
                             
            4'd15: padrao <= {8'b00010000,
                              8'b00110000,
                              8'b00000100,
                              8'b00000100,
                              8'b11000000,
                              8'b11000000,
                              8'b00010000,
                              8'b00001000}; //4
            default: padrao <={8'b11_00_00_11,
                          8'b11_01_01_11,
                          8'b11_11_11_11,
                          8'b11_00_00_11,
                          8'b11_11_11_11,
                          8'b11_00_00_11,
                          8'b11_10_11_11,
                          8'b11_00_00_11};
        endcase
    end

endmodule